.title KiCad schematic
SW1 0 out SW_SPST
V1 Net-_R1-Pad1_ 0 dc 3.3 ac 0
C1 out 0 33p
R1 Net-_R1-Pad1_ out 100k
.control
.tran 2us 100ms 0
.tran 2us 100ms 0
plot d(out)
plot d(out)
.endc
.end
